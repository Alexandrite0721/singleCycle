module InstructionMemory(
	input      [32 -1:0] Address, 
	output reg [32 -1:0] Instruction
);
	
	always @(*)
		case (Address[10:2])
9'd000: Instruction <= 32'h20100000;
9'd001: Instruction <= 32'h20120000;
9'd002: Instruction <= 32'h8e110000;
9'd003: Instruction <= 32'h22230000;
9'd004: Instruction <= 32'h22080004;
9'd005: Instruction <= 32'h22290000;
9'd006: Instruction <= 32'h200a0001;
9'd007: Instruction <= 32'h112a0022;
9'd008: Instruction <= 32'h214cffff;
9'd009: Instruction <= 32'h000a6880;
9'd010: Instruction <= 32'h010d7020;
9'd011: Instruction <= 32'h8dce0000;
9'd012: Instruction <= 32'h0180082a;
9'd013: Instruction <= 32'h14200008;
9'd014: Instruction <= 32'h22520001;
9'd015: Instruction <= 32'h000c6880;
9'd016: Instruction <= 32'h010d7820;
9'd017: Instruction <= 32'h8def0000;
9'd018: Instruction <= 32'h01cf082a;
9'd019: Instruction <= 32'h10200002;
9'd020: Instruction <= 32'h218cffff;
9'd021: Instruction <= 32'h0810000c;
9'd022: Instruction <= 32'h21820001;
9'd023: Instruction <= 32'h214cffff;
9'd024: Instruction <= 32'h000a6880;
9'd025: Instruction <= 32'h010d7020;
9'd026: Instruction <= 32'h8dce0000;
9'd027: Instruction <= 32'h204f0000;
9'd028: Instruction <= 32'h018f082a;
9'd029: Instruction <= 32'h14200007;
9'd030: Instruction <= 32'h000c6880;
9'd031: Instruction <= 32'h010dc020;
9'd032: Instruction <= 32'h8f140000;
9'd033: Instruction <= 32'h23190004;
9'd034: Instruction <= 32'haf340000;
9'd035: Instruction <= 32'h218cffff;
9'd036: Instruction <= 32'h0810001c;
9'd037: Instruction <= 32'h000f7880;
9'd038: Instruction <= 32'h010fc820;
9'd039: Instruction <= 32'haf2e0000;
9'd040: Instruction <= 32'h214a0001;
9'd041: Instruction <= 32'h08100007;
9'd042: Instruction <= 32'hae120000;
9'd043: Instruction <= 32'h20130000;
9'd044: Instruction <= 32'h20080004;
9'd045: Instruction <= 32'h201b07d0;
9'd046: Instruction <= 32'h200f0384;
9'd047: Instruction <= 32'h20180000;
9'd048: Instruction <= 32'h20044000;
9'd049: Instruction <= 32'h20060001;
9'd050: Instruction <= 32'h8d090000;
9'd051: Instruction <= 32'h3122000f;
9'd052: Instruction <= 32'h08100066;
9'd053: Instruction <= 32'h20170100;
9'd054: Instruction <= 32'h00571025;
9'd055: Instruction <= 32'hac820000;
9'd056: Instruction <= 32'h201a0000;
9'd057: Instruction <= 32'h235a0001;
9'd058: Instruction <= 32'h135b0001;
9'd059: Instruction <= 32'h08100039;
9'd060: Instruction <= 32'h8d090000;
9'd061: Instruction <= 32'h00091102;
9'd062: Instruction <= 32'h3042000f;
9'd063: Instruction <= 32'h20c60001;
9'd064: Instruction <= 32'h08100066;
9'd065: Instruction <= 32'h20170200;
9'd066: Instruction <= 32'h00571025;
9'd067: Instruction <= 32'hac820000;
9'd068: Instruction <= 32'h201a0000;
9'd069: Instruction <= 32'h235a0001;
9'd070: Instruction <= 32'h135b0001;
9'd071: Instruction <= 32'h08100045;
9'd072: Instruction <= 32'h8d090000;
9'd073: Instruction <= 32'h00091202;
9'd074: Instruction <= 32'h3042000f;
9'd075: Instruction <= 32'h20c60001;
9'd076: Instruction <= 32'h08100066;
9'd077: Instruction <= 32'h20170400;
9'd078: Instruction <= 32'h00571025;
9'd079: Instruction <= 32'hac820000;
9'd080: Instruction <= 32'h201a0000;
9'd081: Instruction <= 32'h235a0001;
9'd082: Instruction <= 32'h135b0001;
9'd083: Instruction <= 32'h08100051;
9'd084: Instruction <= 32'h8d090000;
9'd085: Instruction <= 32'h00091302;
9'd086: Instruction <= 32'h3042000f;
9'd087: Instruction <= 32'h20c60001;
9'd088: Instruction <= 32'h08100066;
9'd089: Instruction <= 32'h20170800;
9'd090: Instruction <= 32'h00571025;
9'd091: Instruction <= 32'hac820000;
9'd092: Instruction <= 32'h201a0000;
9'd093: Instruction <= 32'h235a0001;
9'd094: Instruction <= 32'h135b0001;
9'd095: Instruction <= 32'h0810005d;
9'd096: Instruction <= 32'h23180001;
9'd097: Instruction <= 32'h170fffce;
9'd098: Instruction <= 32'h22730001;
9'd099: Instruction <= 32'h21080004;
9'd100: Instruction <= 32'h12630049;
9'd101: Instruction <= 32'h0810002e;
9'd102: Instruction <= 32'h20050000;
9'd103: Instruction <= 32'h1045001e;
9'd104: Instruction <= 32'h20a50001;
9'd105: Instruction <= 32'h1045001e;
9'd106: Instruction <= 32'h20a50001;
9'd107: Instruction <= 32'h1045001e;
9'd108: Instruction <= 32'h20a50001;
9'd109: Instruction <= 32'h1045001e;
9'd110: Instruction <= 32'h20a50001;
9'd111: Instruction <= 32'h1045001e;
9'd112: Instruction <= 32'h20a50001;
9'd113: Instruction <= 32'h1045001e;
9'd114: Instruction <= 32'h20a50001;
9'd115: Instruction <= 32'h1045001e;
9'd116: Instruction <= 32'h20a50001;
9'd117: Instruction <= 32'h1045001e;
9'd118: Instruction <= 32'h20a50001;
9'd119: Instruction <= 32'h1045001e;
9'd120: Instruction <= 32'h20a50001;
9'd121: Instruction <= 32'h1045001e;
9'd122: Instruction <= 32'h20a50001;
9'd123: Instruction <= 32'h1045001e;
9'd124: Instruction <= 32'h20a50001;
9'd125: Instruction <= 32'h1045001e;
9'd126: Instruction <= 32'h20a50001;
9'd127: Instruction <= 32'h1045001e;
9'd128: Instruction <= 32'h20a50001;
9'd129: Instruction <= 32'h1045001e;
9'd130: Instruction <= 32'h20a50001;
9'd131: Instruction <= 32'h1045001e;
9'd132: Instruction <= 32'h20a50001;
9'd133: Instruction <= 32'h1045001e;
9'd134: Instruction <= 32'h2002003f;
9'd135: Instruction <= 32'h081000a6;
9'd136: Instruction <= 32'h20020006;
9'd137: Instruction <= 32'h081000a6;
9'd138: Instruction <= 32'h2002005b;
9'd139: Instruction <= 32'h081000a6;
9'd140: Instruction <= 32'h2002004f;
9'd141: Instruction <= 32'h081000a6;
9'd142: Instruction <= 32'h20020066;
9'd143: Instruction <= 32'h081000a6;
9'd144: Instruction <= 32'h2002006d;
9'd145: Instruction <= 32'h081000a6;
9'd146: Instruction <= 32'h2002007d;
9'd147: Instruction <= 32'h081000a6;
9'd148: Instruction <= 32'h20020007;
9'd149: Instruction <= 32'h081000a6;
9'd150: Instruction <= 32'h2002007f;
9'd151: Instruction <= 32'h081000a6;
9'd152: Instruction <= 32'h2002006f;
9'd153: Instruction <= 32'h081000a6;
9'd154: Instruction <= 32'h20020077;
9'd155: Instruction <= 32'h081000a6;
9'd156: Instruction <= 32'h2002007c;
9'd157: Instruction <= 32'h081000a6;
9'd158: Instruction <= 32'h20020058;
9'd159: Instruction <= 32'h081000a6;
9'd160: Instruction <= 32'h2002005e;
9'd161: Instruction <= 32'h081000a6;
9'd162: Instruction <= 32'h20020079;
9'd163: Instruction <= 32'h081000a6;
9'd164: Instruction <= 32'h20020071;
9'd165: Instruction <= 32'h081000a6;
9'd166: Instruction <= 32'h20190001;
9'd167: Instruction <= 32'h10d9ff8d;
9'd168: Instruction <= 32'h23390001;
9'd169: Instruction <= 32'h10d9ff97;
9'd170: Instruction <= 32'h23390001;
9'd171: Instruction <= 32'h10d9ffa1;
9'd172: Instruction <= 32'h23390001;
9'd173: Instruction <= 32'h10d9ffab;
9'd174: Instruction <= 32'h20080f71;
9'd175: Instruction <= 32'hac880000;
9'd176: Instruction <= 32'h081000ae;

			default: Instruction <= 32'h00000000;
		endcase
		
endmodule
